localparam A_WR_SUB					= 76;
localparam PC_WR_JOYPAD_INT		= 75;
localparam PC_WR_SERIAL_INT		= 74;
localparam PC_WR_TIMER_INT			= 73;
localparam PC_WR_LCD_STAT_INT		= 72;
localparam PC_WR_V_BLANK_INT		= 71;
localparam IME_SET					= 70;
localparam IME_RESET					= 69;
localparam A_WR_OR					= 68;
localparam A_WR_AND					= 67;
localparam B_DEC						= 66;
localparam D_DEC						= 65;
localparam A_WR_RRCA					= 64;
localparam A_WR_RLCA					= 63;
localparam A_WR_RRA					= 62;
localparam A_WR_RLA					= 61;
localparam BIT_OP_MSB				= 60;
localparam BIT_OP_LSB				= 58;
localparam CB_IR_WR					= 57;
localparam SP_INC						= 56;
localparam C_DEC						= 55;
localparam A_WR_CPL					= 54;
localparam A_WR_XOR					= 53;
localparam PC_WR_WZ					= 52;
localparam SP_DEC						= 51;
localparam PC_WR_MSB					= 50;
localparam PC_WR_LSB					= 49;
localparam A_INC						= 48;
localparam L_INC						= 47;
localparam H_INC						= 46;
localparam E_INC						= 45;
localparam D_INC						= 44;
localparam C_INC						= 43;
localparam B_INC						= 42;
localparam ADDR_BUS_DEC_WR 		= 41;
localparam ADDR_BUS_INC_WR 		= 40;
localparam ALU_MUX1_MSB				= 39;
localparam ALU_MUX1_LSB				= 36;
localparam ALU_MUX0_MSB				= 35;
localparam ALU_MUX0_LSB				= 32;
localparam ALU_OUT_WR				= 31;
localparam ALU_CNTL_MSB				= 30;
localparam ALU_CNTL_LSB				= 26;
localparam PC_WR						= 25;
localparam SP_WR_MSB					= 24;
localparam SP_WR_LSB					= 23;
localparam MEM_WR						= 22;
localparam A_WR						= 21;
localparam B_WR						= 20;
localparam C_WR						= 19;
localparam D_WR						= 18;
localparam E_WR						= 17;
localparam F_WR						= 16;
localparam H_WR						= 15;
localparam L_WR						= 14;
localparam W_WR						= 13;
localparam Z_WR						= 12;
localparam TMP_WR						= 11;
localparam IR_WR						= 10;
localparam ADDR_BUS_WR				= 9;
localparam PC_INC						= 8;
localparam DATA_BUS_MSB 			= 7;
localparam DATA_BUS_LSB 			= 4;
localparam ADDR_BUS_MSB 			= 3;
localparam ADDR_BUS_LSB 			= 0;

localparam CTRL_MSB					= 76;